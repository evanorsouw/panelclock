library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity linear2logarithmic is
    port (
        lin:	in  std_logic_vector(7 downto 0);
        log:	out std_logic_vector(7 downto 0)
    );
end entity;

architecture linear2logarithmic_arch of linear2logarithmic is
begin
	process (lin) is
	begin 
		case lin is
		when "00000000" => log <= "00000000";
		when "00000001" => log <= "00000000";
		when "00000010" => log <= "00000000";
		when "00000011" => log <= "00000000";
		when "00000100" => log <= "00000000";
		when "00000101" => log <= "00000000";
		when "00000110" => log <= "00000000";
		when "00000111" => log <= "00000000";
		when "00001000" => log <= "00000000";
		when "00001001" => log <= "00000000";
		when "00001010" => log <= "00000000";
		when "00001011" => log <= "00000001";
		when "00001100" => log <= "00000001";
		when "00001101" => log <= "00000001";
		when "00001110" => log <= "00000001";
		when "00001111" => log <= "00000001";
		when "00010000" => log <= "00000001";
		when "00010001" => log <= "00000001";
		when "00010010" => log <= "00000001";
		when "00010011" => log <= "00000001";
		when "00010100" => log <= "00000001";
		when "00010101" => log <= "00000001";
		when "00010110" => log <= "00000010";
		when "00010111" => log <= "00000010";
		when "00011000" => log <= "00000010";
		when "00011001" => log <= "00000010";
		when "00011010" => log <= "00000010";
		when "00011011" => log <= "00000010";
		when "00011100" => log <= "00000010";
		when "00011101" => log <= "00000010";
		when "00011110" => log <= "00000010";
		when "00011111" => log <= "00000010";
		when "00100000" => log <= "00000011";
		when "00100001" => log <= "00000011";
		when "00100010" => log <= "00000011";
		when "00100011" => log <= "00000011";
		when "00100100" => log <= "00000011";
		when "00100101" => log <= "00000011";
		when "00100110" => log <= "00000011";
		when "00100111" => log <= "00000011";
		when "00101000" => log <= "00000011";
		when "00101001" => log <= "00000011";
		when "00101010" => log <= "00000100";
		when "00101011" => log <= "00000100";
		when "00101100" => log <= "00000100";
		when "00101101" => log <= "00000100";
		when "00101110" => log <= "00000100";
		when "00101111" => log <= "00000100";
		when "00110000" => log <= "00000100";
		when "00110001" => log <= "00000100";
		when "00110010" => log <= "00000100";
		when "00110011" => log <= "00000101";
		when "00110100" => log <= "00000101";
		when "00110101" => log <= "00000101";
		when "00110110" => log <= "00000101";
		when "00110111" => log <= "00000101";
		when "00111000" => log <= "00000101";
		when "00111001" => log <= "00000101";
		when "00111010" => log <= "00000101";
		when "00111011" => log <= "00000101";
		when "00111100" => log <= "00000110";
		when "00111101" => log <= "00000110";
		when "00111110" => log <= "00000110";
		when "00111111" => log <= "00000110";
		when "01000000" => log <= "00000110";
		when "01000001" => log <= "00000110";
		when "01000010" => log <= "00000110";
		when "01000011" => log <= "00000110";
		when "01000100" => log <= "00000111";
		when "01000101" => log <= "00000111";
		when "01000110" => log <= "00000111";
		when "01000111" => log <= "00000111";
		when "01001000" => log <= "00000111";
		when "01001001" => log <= "00000111";
		when "01001010" => log <= "00000111";
		when "01001011" => log <= "00000111";
		when "01001100" => log <= "00001000";
		when "01001101" => log <= "00001000";
		when "01001110" => log <= "00001000";
		when "01001111" => log <= "00001000";
		when "01010000" => log <= "00001000";
		when "01010001" => log <= "00001000";
		when "01010010" => log <= "00001000";
		when "01010011" => log <= "00001000";
		when "01010100" => log <= "00001001";
		when "01010101" => log <= "00001001";
		when "01010110" => log <= "00001001";
		when "01010111" => log <= "00001001";
		when "01011000" => log <= "00001001";
		when "01011001" => log <= "00001001";
		when "01011010" => log <= "00001001";
		when "01011011" => log <= "00001010";
		when "01011100" => log <= "00001010";
		when "01011101" => log <= "00001010";
		when "01011110" => log <= "00001010";
		when "01011111" => log <= "00001010";
		when "01100000" => log <= "00001010";
		when "01100001" => log <= "00001010";
		when "01100010" => log <= "00001011";
		when "01100011" => log <= "00001011";
		when "01100100" => log <= "00001011";
		when "01100101" => log <= "00001011";
		when "01100110" => log <= "00001011";
		when "01100111" => log <= "00001011";
		when "01101000" => log <= "00001011";
		when "01101001" => log <= "00001100";
		when "01101010" => log <= "00001100";
		when "01101011" => log <= "00001100";
		when "01101100" => log <= "00001100";
		when "01101101" => log <= "00001100";
		when "01101110" => log <= "00001100";
		when "01101111" => log <= "00001101";
		when "01110000" => log <= "00001101";
		when "01110001" => log <= "00001101";
		when "01110010" => log <= "00001101";
		when "01110011" => log <= "00001101";
		when "01110100" => log <= "00001101";
		when "01110101" => log <= "00001101";
		when "01110110" => log <= "00001110";
		when "01110111" => log <= "00001110";
		when "01111000" => log <= "00001110";
		when "01111001" => log <= "00001110";
		when "01111010" => log <= "00001110";
		when "01111011" => log <= "00001110";
		when "01111100" => log <= "00001111";
		when "01111101" => log <= "00001111";
		when "01111110" => log <= "00001111";
		when "01111111" => log <= "00001111";
		when "10000000" => log <= "00001111";
		when "10000001" => log <= "00010000";
		when "10000010" => log <= "00010000";
		when "10000011" => log <= "00010000";
		when "10000100" => log <= "00010000";
		when "10000101" => log <= "00010000";
		when "10000110" => log <= "00010000";
		when "10000111" => log <= "00010001";
		when "10001000" => log <= "00010001";
		when "10001001" => log <= "00010001";
		when "10001010" => log <= "00010001";
		when "10001011" => log <= "00010001";
		when "10001100" => log <= "00010010";
		when "10001101" => log <= "00010010";
		when "10001110" => log <= "00010010";
		when "10001111" => log <= "00010010";
		when "10010000" => log <= "00010010";
		when "10010001" => log <= "00010011";
		when "10010010" => log <= "00010011";
		when "10010011" => log <= "00010011";
		when "10010100" => log <= "00010011";
		when "10010101" => log <= "00010011";
		when "10010110" => log <= "00010100";
		when "10010111" => log <= "00010100";
		when "10011000" => log <= "00010100";
		when "10011001" => log <= "00010100";
		when "10011010" => log <= "00010101";
		when "10011011" => log <= "00010101";
		when "10011100" => log <= "00010101";
		when "10011101" => log <= "00010101";
		when "10011110" => log <= "00010101";
		when "10011111" => log <= "00010110";
		when "10100000" => log <= "00010110";
		when "10100001" => log <= "00010110";
		when "10100010" => log <= "00010110";
		when "10100011" => log <= "00010111";
		when "10100100" => log <= "00010111";
		when "10100101" => log <= "00010111";
		when "10100110" => log <= "00010111";
		when "10100111" => log <= "00011000";
		when "10101000" => log <= "00011000";
		when "10101001" => log <= "00011000";
		when "10101010" => log <= "00011000";
		when "10101011" => log <= "00011001";
		when "10101100" => log <= "00011001";
		when "10101101" => log <= "00011001";
		when "10101110" => log <= "00011010";
		when "10101111" => log <= "00011010";
		when "10110000" => log <= "00011010";
		when "10110001" => log <= "00011010";
		when "10110010" => log <= "00011011";
		when "10110011" => log <= "00011011";
		when "10110100" => log <= "00011011";
		when "10110101" => log <= "00011100";
		when "10110110" => log <= "00011100";
		when "10110111" => log <= "00011100";
		when "10111000" => log <= "00011101";
		when "10111001" => log <= "00011101";
		when "10111010" => log <= "00011101";
		when "10111011" => log <= "00011110";
		when "10111100" => log <= "00011110";
		when "10111101" => log <= "00011110";
		when "10111110" => log <= "00011111";
		when "10111111" => log <= "00011111";
		when "11000000" => log <= "00011111";
		when "11000001" => log <= "00100000";
		when "11000010" => log <= "00100000";
		when "11000011" => log <= "00100000";
		when "11000100" => log <= "00100001";
		when "11000101" => log <= "00100001";
		when "11000110" => log <= "00100010";
		when "11000111" => log <= "00100010";
		when "11001000" => log <= "00100010";
		when "11001001" => log <= "00100011";
		when "11001010" => log <= "00100011";
		when "11001011" => log <= "00100100";
		when "11001100" => log <= "00100100";
		when "11001101" => log <= "00100100";
		when "11001110" => log <= "00100101";
		when "11001111" => log <= "00100101";
		when "11010000" => log <= "00100110";
		when "11010001" => log <= "00100110";
		when "11010010" => log <= "00100111";
		when "11010011" => log <= "00100111";
		when "11010100" => log <= "00101000";
		when "11010101" => log <= "00101000";
		when "11010110" => log <= "00101001";
		when "11010111" => log <= "00101001";
		when "11011000" => log <= "00101010";
		when "11011001" => log <= "00101011";
		when "11011010" => log <= "00101011";
		when "11011011" => log <= "00101100";
		when "11011100" => log <= "00101100";
		when "11011101" => log <= "00101101";
		when "11011110" => log <= "00101110";
		when "11011111" => log <= "00101110";
		when "11100000" => log <= "00101111";
		when "11100001" => log <= "00110000";
		when "11100010" => log <= "00110001";
		when "11100011" => log <= "00110001";
		when "11100100" => log <= "00110010";
		when "11100101" => log <= "00110011";
		when "11100110" => log <= "00110100";
		when "11100111" => log <= "00110101";
		when "11101000" => log <= "00110110";
		when "11101001" => log <= "00110111";
		when "11101010" => log <= "00111000";
		when "11101011" => log <= "00111001";
		when "11101100" => log <= "00111010";
		when "11101101" => log <= "00111011";
		when "11101110" => log <= "00111100";
		when "11101111" => log <= "00111110";
		when "11110000" => log <= "00111111";
		when "11110001" => log <= "01000000";
		when "11110010" => log <= "01000010";
		when "11110011" => log <= "01000100";
		when "11110100" => log <= "01000110";
		when "11110101" => log <= "01001000";
		when "11110110" => log <= "01001010";
		when "11110111" => log <= "01001100";
		when "11111000" => log <= "01001111";
		when "11111001" => log <= "01010010";
		when "11111010" => log <= "01010101";
		when "11111011" => log <= "01011010";
		when "11111100" => log <= "01011111";
		when "11111101" => log <= "01100101";
		when "11111110" => log <= "01101111";
		when "11111111" => log <= "01111111";
		end case;
	end process;
end architecture;
